module full_adder(	input [1:0] a,
			input [1:0] b, 
			input [1:0] c_in,
			output [1:0] sum,
			output [1:0] c_out
);




endmodule

